module adder_32 (
    input[31:0] in1, in2,
    output[31:0] out
);
    out = in1 + in2;
    
endmodule