module registers (
    input[31:0] data_in, wr_idx, r1_idx, r2_idx,
    input wr_en, reset, clk,
    output[31:0] reg_1, data_2
);
    


endmodule