module full_system (

    
endmodule